library verilog;
use verilog.vl_types.all;
entity dec_imp_tb is
end dec_imp_tb;
