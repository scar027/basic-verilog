module xor_gate(y,a,b);
  input a, b;
  output y;
  xor xor1(y,a,b);
endmodule  