module nor_gate(y,a,b);
  input a, b;
  output y;
  nor no1(y,a,b);
endmodule  
