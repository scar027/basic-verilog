module not_gate(y,a);
  input a;
  output y;
  not n1(y,a);
endmodule