library verilog;
use verilog.vl_types.all;
entity sr_latch_nor_tb is
end sr_latch_nor_tb;
