module and_gate(y,a,b);
  input a, b;
  output y;
  and a1(y,a,b);
endmodule  
