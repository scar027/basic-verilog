library verilog;
use verilog.vl_types.all;
entity rca_test is
end rca_test;
