library verilog;
use verilog.vl_types.all;
entity fulladder_test is
end fulladder_test;
