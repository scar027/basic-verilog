module decoder_implementation (x, y, y0, y1, y2, y3, y4, 
y5, y6, y7, y8, y9, y10, 
y11, y12, y13, y14, y15, a, b, c, d);
  input a, b, c, d;
  output x, y, y0, y1, y2, y3, y4, y5, 
  y6, y7, y8, y9, y10, y11, y12, y13, y14, y15;
  reg x, y, y0, y1, y2, y3, y4, y5, 
  y6, y7, y8, y9, y10, y11, y12, y13, y14, y15;
  always @ (a or b or c or d)
  begin
    case({a,b,c,d})
      4'b0000 : begin y0 = 1; y1 = 0; y2 = 0; 
      y3 = 0 ; y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; 
      y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0001 : begin y0 = 0; y1 = 1; y2 = 0; 
      y3 = 0; y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0010 : begin y0 = 0; y1 = 0; y2 = 1; y3 = 0; 
      y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0011 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 1
      y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0100 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0 ;
       y4 = 1; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; 
      y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0101 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0; 
      y4 = 0; y5 = 1; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; 
      y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0110 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0;
       y4 = 0; y5 = 0; 
                      
      y6 = 1; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b0111 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0;
      y4 = 0; y5 = 0; 
      y6 = 0; y7 = 1; y8 = 0; y9 = 0; 
      y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b1000 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0; 
      y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 1; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b1001 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0; 
      y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 1; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b1010 : begin y0 = 0; y1 = 0; y2 = 0; 
      y3 = 0; y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 1; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b1011 : begin y0 = 0; y1 = 0; y2 = 0;
      y3 = 0; y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; 
      y9 = 0; y10 = 0; y11 = 1; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 0; end
      4'b1100 : begin y0 = 0; y1 = 0; y2 = 0; 
      y3 = 0; y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 1; y13 = 0; y14 = 0; y15 = 0; end
      4'b1101 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0; 
      y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 1; y14 = 0; y15 = 0; end
      4'b1110 : begin y0 = 0; y1 = 0; y2 = 0; y3 = 0;
       y4 = 0; y5 = 0; 
       y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 1; y15 = 0; end
      4'b1111 : begin y0 = 0; y1 = 0; y2 = 0; 
      y3 = 0; y4 = 0; y5 = 0; 
      y6 = 0; y7 = 0; y8 = 0; y9 = 0; y10 = 0; y11 = 0; 
      y12 = 0; y13 = 0; y14 = 0; y15 = 1; end                                                                                                                                
      
    endcase
    
    assign x = (y2|y3|y10|y11|y12|y13|y14|y15);
    assign y = (y4|y6|y7|y8|y10|y11|y12|y14|y15);
    
  end
endmodule        
