library verilog;
use verilog.vl_types.all;
entity decoder_implementation is
    port(
        x               : out    vl_logic;
        y               : out    vl_logic;
        y0              : out    vl_logic;
        y1              : out    vl_logic;
        y2              : out    vl_logic;
        y3              : out    vl_logic;
        y4              : out    vl_logic;
        y5              : out    vl_logic;
        y6              : out    vl_logic;
        y7              : out    vl_logic;
        y8              : out    vl_logic;
        y9              : out    vl_logic;
        y10             : out    vl_logic;
        y11             : out    vl_logic;
        y12             : out    vl_logic;
        y13             : out    vl_logic;
        y14             : out    vl_logic;
        y15             : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic
    );
end decoder_implementation;
