library verilog;
use verilog.vl_types.all;
entity mux_41_case is
    port(
        \out\           : out    vl_logic;
        i0              : in     vl_logic;
        i1              : in     vl_logic;
        i2              : in     vl_logic;
        i3              : in     vl_logic;
        s1              : in     vl_logic;
        s0              : in     vl_logic
    );
end mux_41_case;
