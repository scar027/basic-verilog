library verilog;
use verilog.vl_types.all;
entity mux_41_tb is
end mux_41_tb;
