library verilog;
use verilog.vl_types.all;
entity ckt_tb is
end ckt_tb;
