library verilog;
use verilog.vl_types.all;
entity demuxtest is
end demuxtest;
