library verilog;
use verilog.vl_types.all;
entity beh_cond_tb is
end beh_cond_tb;
