library verilog;
use verilog.vl_types.all;
entity halfadder_test is
end halfadder_test;
