module nand_gate(y,a,b);
  input a, b;
  output y;
  nand nal(y,a,b);
endmodule  

