module or_gate(y,a,b);
  input a, b;
  output y;
  or o1(y,a,b);
endmodule  