library verilog;
use verilog.vl_types.all;
entity halfadderiftb is
end halfadderiftb;
