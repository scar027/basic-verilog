library verilog;
use verilog.vl_types.all;
entity decoder_21_tb is
end decoder_21_tb;
